/* 
    This is just the kogge-stone adder written for VLSI ported to system verilog
 */

 module 4bit_ksadd;

    wire 

 endmodule;