module and(in 1, )